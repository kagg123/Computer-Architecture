`timescale 1ns/10ps
module cpu(input logic clk, reset);
	
	logic [31:0] instruction;
	logic [31:0] instructionOut;
	logic        zeroFlag, zero_cbzcheck, reg2Loc, unCondBr, isBL, isCbz, isBlt,
	             negFlag, overflowFlag, carry_outFlag;
	logic [1:0]  brTaken;
	logic [4:0] Rd [3:0];
	logic [4:0] Rm, Rn;
	//logic [4:0] RdOut, RmOut, RnOut;
	logic [8:0] Imm9;
	logic [11:0] Imm12;
	logic [18:0] condAddr19;
	logic [25:0] condAddr26;
	logic [63:0] forwardCtrlOneOutput, pc_output;
	
	// instantiate the dataPath module
	
	logic [1:0] forwardCtrlOne ;
	logic [1:0] forwardCtrlTwo;
	logic [3:0] regWrite;
	logic [2:0] memWrite;
	logic [1:0] flagEn;
	
	logic [1:0] aluSrc;
	logic [2:0] aluOp [1:0];
	logic [1:0] memToReg [2:0];
	// logic Rd1, Rd2; 

	// paramDFF #(parameter WIDTH = 5) pdff1 (.d(RdOut), .q(Rd1), .reset, .clk);
	// paramDFF #(parameter WIDTH = 5) pdff2 (.d(Rd1), .q(Rd2)), .reset, .clk);
	forwardingUnit fd (.Rd1(Rd[2]), .Rd2(Rd[1]), .Rm, .Rn, .forwardCtrlOne, .forwardCtrlTwo, .regWrite1(regWrite[2]), .regWrite2(regWrite[1]));
	
	
	//control path registers
	IFID r1 (.instruction(instruction), .zeroFlag, .negFlag(negFlag), .overflowFlag(overflowFlag), .clk, .reset, .Rd(Rd[3]), .Rm, .Rn,
			.Imm12, .Imm9, .condAddr19, .condAddr26, .brTaken, .aluSrc, .memToReg(memToReg[2]), .aluOp(aluOp[1]),
			.reg2Loc, .memWrite(memWrite[2]), .regWrite(regWrite[3]), .unCondBr, .flagEn(flagEn[1]), .isCbz, .isBlt);

	IDEX r2(.clk, .reset, .aluOp(aluOp[1]), .memToReg(memToReg[2]), .memWrite(memWrite[2]), .regWrite(regWrite[3]), .flagEn(flagEn[1]), 
			 .Rd(Rd[3]), .RdOut(Rd[2]),  .aluOpOut(aluOp[0]), .memToRegOut(memToReg[1]), .memWriteOut(memWrite[1]), 
			 .regWriteOut(regWrite[2]), .flagEnOut(flagEn[0]));
	
    EXMEM r3 (.clk, .reset, .memToReg(memToReg[1]), .memWrite(memWrite[1]), .regWrite(regWrite[2]), .Rd(Rd[2]), 
				.RdOut(Rd[1]), .memToRegOut(memToReg[0]), .memWriteOut(memWrite[0]), .regWriteOut(regWrite[1]));
	
	MEMWR r4 (.clk, .reset, .regWrite(regWrite[1]),  .Rd(Rd[1]), .RdOut(Rd[0]), .regWriteOut(regWrite[0]));
	
	
	//dataPath IFID Regsiter
	paramDFF #(.WIDTH(32)) ifidDataRegister (.d(instruction), .q(instructionOut), .reset, .clk);

	logic [1:0] brTakenActual;
	logic [1:0] brTakenisCbzBlt [2:0];
	logic xorOverflowNegative;

	xor #0.05 x1 (xorOverflowNegative, negFlag, overflowFlag);

	assign brTakenisCbzBlt[2] = {1'b0, xorOverflowNegative};
	assign brTakenisCbzBlt[1] = {1'b0, zero_cbzcheck};
	assign brTakenisCbzBlt[0] = brTaken;

	mux2x3_1 m9000 (.muxOutput(brTakenActual), .muxInputs(brTakenisCbzBlt), .select({isBlt, isCbz}));
	
	instructfetch fetch (.reset, .clk, .uncondBr(unCondBr), .brTaken(brTakenActual), .condAddr19, 
	                     .condAddr26, .forwardCtrlOneOutput, .instruction, .pc_output);
								
	dataPath path (.reg2Loc, .regWrite(regWrite[0]), .clk, .memWrite(memWrite[0]), .flagEn(flagEn[0]), .reset, 
                  .aluSrc(aluSrc), .memToReg(memToReg[0]), .aluOp(aluOp[0]), .forwardCtrlOne, .forwardCtrlTwo, 
				  .Rd(Rd[0]), .Rm, .Rn, .Imm9, .Imm12,
				      .pc_output, .negFlag, .zeroFlag, .zero_cbzcheck, .overflowFlag, .carry_outFlag, .forwardCtrlOneOutput);
						
	
endmodule


module cpu_testbench();

	logic clk, reset;
	
	cpu dut (.clk, .reset);
	
	// Set up the clock.   
	parameter CLOCK_PERIOD = 100000;   
	initial begin    
		clk <= 0;    
		forever #( CLOCK_PERIOD / 2 ) clk <= ~clk;   
	end 
	
	
	initial begin
										@( posedge clk );    
		 reset <= 1'b1;         @( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
		 reset <= 1'b0;			@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
		 reset <= 1'b0;			@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
																				@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk ); 
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );
										@( posedge clk );


										
		 $stop; // End the simulation.
		 
	end
	
	
endmodule




